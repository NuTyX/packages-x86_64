msgid ""
msgstr ""
"Project-Id-Version: NuTyX Configuration tool\n"
"PO-Revision-Date: 2014-08-07+2000\n"
"Last-Translator: https://translate.google.se/#fr/sv/\n"
"Language-Team: Swedish\n"
"Language: sv \n"
"MIME-Version: 1.0\n"
"Content-Type: text/plain; charset=UTF-8\n"
"Content-Transfer-Encoding: 8bit\n"

msgid "Settings"
msgstr "Inställningar"

msgid "Keyboard Layout"
msgstr "Tangentbordslayout"

msgid "Choose available"
msgstr "Välj tillgängliga"

msgid "ERROR configuration"
msgstr "Konfigurationsfel"

msgid "Please try again"
msgstr "Försök igen"

msgid "Network card"
msgstr "Nätverkskort"

msgid "Select the card"
msgstr "Välj kort"

msgid "Card to configure"
msgstr "Kort att konfigurera"

msgid "Configuration of"
msgstr "Konfiguration av"

msgid "Configuration mode"
msgstr "Konfigurationsläge"

msgid "Auto"
msgstr "Auto"

msgid "Man"
msgstr "Man"

msgid "IP address automatically set from DHCP server"
msgstr "IP adress häntas automatiskt från DHCP-servern"

msgid "Manually specify parameters"
msgstr "Ange parametrar manuellt"

msgid "Enter an IP address"
msgstr "Ange en IP-adress"

msgid "Enter a broadcast address"
msgstr "Ange en broadcast-adress"

msgid "in most cases the current value can be used"
msgstr "i de flesta fall kan det aktuella värdet kan användas"

msgid "Enter the subnet mask"
msgstr "Ange nätmasken"

msgid "Enter the gateway address"
msgstr "Ange gateway-adress"

msgid "it is normally the address of your router access point"
msgstr "det är normalt adressen för din router åtkomstpunkt"

msgid "Enter the DNS address"
msgstr "Ange DNS-adress"

msgid "DNS Search Suffix"
msgstr "DNS-sökning Suffix"

msgid "Enter the domain name"
msgstr "Ange domännamn"

msgid "this is only need if you are in a subdomain"
msgstr "detta behövs bara om du är i en underdomän"

msgid "Most of the time it's not need"
msgstr "Men oftast behövs det inte göras"

msgid "Start the service"
msgstr "Starta tjänsten"

msgid "Checking the configuration, returning true or false"
msgstr "Analyserar inställningar, returnerar sant eller falskt"

msgid "Show the network configuration"
msgstr "Visa nätverkskonfigurationen"

msgid "Show the keyboard configuration"
msgstr "Visa tangentbordskonfigurationen"

msgid "Show the date and time settings"
msgstr "Visa tids och datum inställningar"

msgid "Show the timezone and time adjustment"
msgstr "Visa tids zon och tid inställningar"

msgid "Show all configurations"
msgstr "Visa all konfiguration"

msgid "Configure the language"
msgstr "Språk inställning"

msgid "Configure the keyboard"
msgstr "Konfigurera tangentbordet"

msgid "Configure the network"
msgstr "Konfigurera nätverket"

msgid "Date and time settings"
msgstr "Datum och tid inställningar"

msgid "Add a user to the system"
msgstr "Lägg till en användare i systemet"

msgid "Configure the system"
msgstr "Konfigurera systemet"

msgid "Install NuTyX"
msgstr "Installera NuTyX"

msgid "Use the arrows keys to change the values"
msgstr "Använd piltangenterna för att ändra värdena"

msgid "Coordinated Universal Time or Local Time ?"
msgstr "Coordinated Universal Time eller Lokal tid ?"

msgid "The hardware clock is set to"
msgstr "Maskinvaruklockan är inställd på"

msgid "Do you want to use this time as Coordinated Universal Time ?"
msgstr "Vill du använda denna tid som Coordinated Universal Time ?"

msgid "so that the summer/winter time is changed automatically"
msgstr "så att sommar / vintertid ändras automatiskt"

msgid "Please enter the date"
msgstr "Vänligen ange datum"

msgid "Please enter the time"
msgstr "Ange tiden"

msgid "Configuration of the boot of the computer (GRUB)"
msgstr "Konfiguration av boot inställingar av datorn (GRUB)"

msgid "Select the disk on which you want to modify the MBR"
msgstr "Välj den disk som du vill ändra MBR på"

msgid "Select the partition on which you want to place the GRUB files"
msgstr "Välj den partition som vill placera GRUB-filerna på"

msgid "Note that the destination partition can contain NuTyX or any other distribution"
msgstr "Observera att destinationen partition kan innehålla NuTyX eller någon annan distribution"

msgid "No boot process configured"
msgstr "Ingen boot process konfigurerad"

msgid "You have installed NuTyX without configuring the boot process"
msgstr "Du har installerat NuTyX utan konfiguration av boot process"

msgid "Are you sure, you want to cancel the process ?"
msgstr "Är du säker på att du vill avbryta processen ?"

msgid "You already have a copy of the original MBR, I will not make a backup of it"
msgstr "Du har redan en kopia av den ursprungliga MBR, jag gör ingen backup på den"

msgid "Everything OK, do you want to modify"
msgstr "Allt är OK, vill du ändra"

msgid "Something went wrong probably the file system is not supported"
msgstr "Något gick fel, förmodligen stöds inte filsystemet"

msgid "A new"
msgstr "En ny"

msgid "has been created"
msgstr "har skapats"

msgid "it has been adapted to launch the Maintenance system of NuTyX"
msgstr "Den är anpassad för att starta underhålls systemet i NuTyX"

msgid "if you choose"
msgstr "Om du väljer"

msgid "an simplify VI editor will allow you to modify it"
msgstr "en förenklad VI editor låter dig ändra den"

msgid "Enter the edit mode"
msgstr "Starta redigeringsläge"

msgid "Exit the edit mode"
msgstr "Avsluta redigeringsläge"

msgid "Cancel the modifications and exit VI"
msgstr "Ångra ändringarna och gå ur VI"

msgid "Save and exit VI"
msgstr "Spara och gå ur VI"

msgid "Good to know"
msgstr "Bra att veta"

msgid "Main Menu"
msgstr "Huvudmeny"

msgid "Welcome to the NuTyX installer"
msgstr "Välkommen till NuTyX installationen"

msgid "Create all your partitions"
msgstr "Skapa alla dina partitioner"

msgid "Format a partition"
msgstr "Formatera en partition"

msgid "Configure the boot of the PC"
msgstr "Konfigurera datorns uppstartsprocess"

msgid "Reboot the PC"
msgstr "Starta om datorn"

msgid "Press OK to reboot the computer"
msgstr "Tryck OK för att starta om datorn"

msgid "optional"
msgstr "valfritt"

msgid "Install"
msgstr "Installera"

msgid "Partitioning"
msgstr "Partitionering"

msgid "Format"
msgstr "Formatering"

msgid "Boot"
msgstr "Boot"

msgid "Keyboard"
msgstr "Tangentbord"

msgid "Network"
msgstr "Nätverk"

msgid "Clock"
msgstr "Klocka"

msgid "Restart"
msgstr "Omstart"

msgid "Yes"
msgstr "Ja"

msgid "Choose the disk you want to use for this operation"
msgstr "Välj hårddisken som du vill använda för denna operation"

msgid "Choose the partition you want to use for this operation"
msgstr "Välj partition som du vill använda för denna operation"

msgid "Available file systems"
msgstr "Tillgängliga filsystem"

msgid "Choose the file system you want to use for the partition"
msgstr "Välj filsystemet som du vill använda för partitionen"

msgid "High performance journaling file system create by SGI"
msgstr "Högprestandafilsystem skapad av SGI"

msgid "Journaling file system create by IBM"
msgstr "Journalförings fil system skapad av IBM"

msgid "Very stable file system but not maintain anymore"
msgstr "Mycket stabilt filsystem som inte upprätthålls längre"

msgid "Next generation of Ext3 file system"
msgstr "Nästa generation av Ext3 filsystemet"

msgid "Journaling version of Ext2 file system"
msgstr "Journalförings version av ext2 filsystem"

msgid "Standard file system Ext2"
msgstr "Standard fil system Ext2"

msgid "New promising file system"
msgstr "Lovande nytt fil system"

msgid "Launch the format process ?"
msgstr "Starta formatierings processen ?"

msgid "The partition"
msgstr "Partitionen"

msgid "will be formatted in"
msgstr "kommer att formateras som"

msgid "Are you sure you want to continue ?"
msgstr "Är du säker på att du vill fortsätta ?"

msgid "No disk available"
msgstr "Ingen hårddisk tillgänglig"

msgid "Please stop the PC and install a harddisk"
msgstr "Stäng datorn och installera en hårddisk"

msgid "No partition available"
msgstr "Ingen partition tillgänglig"

msgid "Please create/modify yours partitions"
msgstr "Skapa / ändra dina partitioner"

msgid "Choose your favorite tool"
msgstr "Välj ditt favorit verktyg"

msgid "Basic partitioning tool"
msgstr "Grundläggande partitioneringsverktyg"

msgid "Advanced partitioning tool"
msgstr "Avancerad partitioneringsverktyg"

msgid "Partitioning of the disk"
msgstr "Partitionering av disken"

msgid "Open a console"
msgstr "Öppna en konsol"

msgid "Please wait"
msgstr "Var god vänta"

msgid "This is a very basic tool, do not expect too much"
msgstr "Detta är ett mycket grundläggande verktyg, förvänta dig inte för mycket"

msgid "It will ask you on which partition you want to install NuTyX"
msgstr "Den kommer att fråga dig om vilken partition du vill installera NuTyX på"

msgid "If not yet created/formatted, it will prompt you to do so"
msgstr "Om den ännu inte är skapad / formaterad, kommer den att fråga dig att göra det"

msgid "No future plan to make this installer more sophisticated"
msgstr "Ingen framtida plan för att göra den här installeraren mer sofistikerade"

msgid "NuTyX goes on"
msgstr "NuTyX läggs på"

msgid "only ONE partition"
msgstr "endast en partition"

msgid "ONE exception, GRUB can be part of it, installed on a separate partition or not installed at all"
msgstr "Ett undantag, GRUB kan vara en del av den, installeras på en separerad partition, eller inte installerad alls"

msgid "As NuTyX users, we recommand you to install GRUB on a separate partition"
msgstr "Som NuTyX användare, rekommenderar vi dig att installera GRUB på en separat partition"

msgid "To do so"
msgstr "För att göra så"

msgid "Install GRUB first, then NuTyX"
msgstr "Installerar GRUB först, sedan NuTyX"

msgid "Have fun"
msgstr "Ha det så kul"

msgid "Thank you for installing NuTyX"
msgstr "Tack för att du installerar NuTyX"

msgid "Help"
msgstr "Hjälp"

msgid "How to do it"
msgstr "Anvisningar"

msgid "A copy of the original MBR is saved in the folder /boot/grub of your NuTyX. It will then be possible to restore it if need"
msgstr "En kopia av original MBR sparas i mappen /boot/grub i din NuTyX. Den kan då återställas om det behövs"

msgid "The name you enter is invalid"
msgstr "Namnet du angav är inte giltigt"

msgid "The name you enter is already register on the system"
msgstr "Namnet du angav är redan upptaget"

msgid "The description you enter is invalid"
msgstr "Beskrivningen du angav är inte giltig"

msgid "Name of the user"
msgstr "Användarnamnet"

msgid "Add a description for the user"
msgstr "Lägg till en användar beskrivning"

msgid "Name or Description of the user"
msgstr "Benämning av användaren"

msgid "Password"
msgstr "Lösenord"

msgid "Enter a new password"
msgstr "Ange ett nytt lösenord"

msgid "Confirm the new password"
msgstr "Bekräfta det nya lösenordet"

msgid "Passwords are differents, please try again"
msgstr "Lösenorden är inte lika, var god försök igen"

msgid "Do you want to try again"
msgstr "Vill du försöka igen?"

msgid "Please run this command as root"
msgstr "Var god kör kommandot som root"

msgid "Sync the HD"
msgstr "Synka HD"

msgid "Emptying memory"
msgstr "Tömmer minnet"

msgid "Swap partition not found"
msgstr "Swap partitionen ej funnen"

msgid "recommended"
msgstr "rekommenderad"

msgid "skilled"
msgstr "erfaren"

msgid "Configure the wireless access point"
msgstr "Konfigurera den tradlösa atkomstpunkten"

msgid "Configuration of a wireless access point for"
msgstr "Konfiguration av den tradlösa atkomstpunkten för"

msgid "Choose the name of the wireless access point"
msgstr "Choose the name of"

msgid "Enter the password of"
msgstr "Enter the password of"

msgid "File"
msgstr "File"

msgid "successfully created"
msgstr "successfully created"

msgid "Cannot create"
msgstr "Cannot create"

msgid "Erase"
msgstr "Erase"

msgid "Configure automatic update"
msgstr "Configure automatic update"

msgid "Would you like to enable automatic update"
msgstr "Would you like to enable automatic update"

msgid "Make shure you reserve the first partition for ESP"
msgstr "Make shure you reserve the first partition for ESP"

msgid "At partitioning, declare the first partition as EFI System"
msgstr "At partitioning, declare the first partition as EFI System"

msgid "EFI partition not found"
msgstr "EFI partition not found"

msgid "GPT partition table not found"
msgstr "GPT partition table not found"

msgid "This installation won't boot again ..."
msgstr "This installation won't boot again ..."

msgid "You can remove the ISO media now."
msgstr "Du kan ta bort media som innehåller ISO nu."

msgid "Advanced Menu"
msgstr "Avancerad meny"

msgid "Advanced"
msgstr "Avancerad"

msgid "Main"
msgstr "Huvud"
